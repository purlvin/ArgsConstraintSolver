
constraint Var_1 { 
  Var1 inside {[10:20]};
}

constraint Var_2 {
  Var2 dist {'h1:=10,'h2:=10};
}

